** sch_path: /home/Joerdson/Downloads/Up_Converter_5GHz.sch
.subckt Mixer5GHz RFN RFP VDC IFP IFN GND ICC LON2 LOP2 VCC2 ICC2 GND2 IDC VCTR2 VCTR VCC
XN6 RFN LON net2 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XRL2 RFN VDC rppd w=4.72e-6 l=8.82e-6 m=1 b=0
XRL1 RFP VDC rppd w=4.72e-6 l=8.82e-6 m=1 b=0
XN8 RFN LOP net3 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XN7 RFP LON net3 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XN5 RFP LOP net2 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XN4 net3 IFN net1 GND sg13_lv_nmos w=160.0u l=0.13u ng=20 m=1
XN3 net2 IFP net1 GND sg13_lv_nmos w=160.0u l=0.13u ng=20 m=1
XN1 IDC IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XN2 net1 IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XN11 LOP LON net4 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XN12 LON LOP net4 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XN9 ICC ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XN10 net4 ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XC1 VCC LOP cap_cmim w=6.62e-6 l=2.42e-6 m=1
XR1 LOP VCC rppd w=10.77e-6 l=8.92e-6 m=1 b=0
XC2 VCC LON cap_cmim w=6.62e-6 l=2.42e-6 m=1
XR2 LON VCC rppd w=10.77e-6 l=8.92e-6 m=1 b=0
XN15 LOP2 LON2 net5 GND2 sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XN16 LON2 LOP2 net5 GND2 sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XN13 ICC2 ICC2 GND2 GND2 sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XN14 net5 ICC2 GND2 GND2 sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XC4 VCC2 LOP2 cap_cmim w=8.73e-6 l=9.42e-6 m=1
XR4 LOP2 VCC2 rppd w=10.77e-6 l=8.92e-6 m=1 b=0
XC5 VCC2 LON2 cap_cmim w=8.73e-6 l=9.42e-6 m=1
XR5 LON2 VCC2 rppd w=10.77e-6 l=8.92e-6 m=1 b=0
L4 VCC2 LOP2 2.006n m=1
L1 VCC LOP 2.006n m=1
L2 VCC LON 2.006n m=1
L5 VCC2 LON2 2.006n m=1
XC6 LOP2 VCTR2 LON2 net5 sg13_hv_svaricap W=9.74e-6 L=0.8e-6 Nx=2
XC3 LOP VCTR LON GND sg13_hv_svaricap W=9.74e-6 L=0.8e-6 Nx=2
XM1 GND net7 net6 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM2 net7 net6 VCC VCC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM3 GND net9 net8 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM4 net9 net8 VCC VCC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM5 GND net11 net10 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM6 net11 net10 VCC VCC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM7 GND net13 net12 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM8 net13 net12 VCTR VCTR sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM9 GND net15 net14 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM10 net15 net14 VCTR VCTR sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM11 GND net17 net16 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM12 net17 net16 VCTR VCTR sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM13 GND net19 net18 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM14 net19 net18 VDC VDC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM15 GND net21 net20 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM16 net21 net20 VDC VDC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM17 GND net23 net22 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM18 net23 net22 VDC VDC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM19 GND net25 net24 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM20 net25 net24 ICC ICC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM21 GND net27 net26 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM22 net27 net26 ICC ICC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM23 GND net29 net28 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM24 net29 net28 ICC ICC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM25 GND net31 net30 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM26 net31 net30 IDC IDC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM27 GND net33 net32 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM28 net33 net32 IDC IDC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM29 GND net35 net34 GND sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM30 net35 net34 IDC IDC sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM31 GND2 net37 net36 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM32 net37 net36 VCTR2 VCTR2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM33 GND2 net39 net38 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM34 net39 net38 VCTR2 VCTR2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM35 GND2 net41 net40 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM36 net41 net40 VCTR2 VCTR2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM37 GND2 net43 net42 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM38 net43 net42 ICC2 ICC2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM39 GND2 net45 net44 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM40 net45 net44 ICC2 ICC2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM41 GND2 net47 net46 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM42 net47 net46 ICC2 ICC2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM49 GND2 net49 net48 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM50 net49 net48 VCC2 VCC2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM51 GND2 net51 net50 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM52 net51 net50 VCC2 VCC2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
XM53 GND2 net53 net52 GND2 sg13_lv_nmos w=250u l=0.13u ng=25 m=1
XM54 net53 net52 VCC2 VCC2 sg13_lv_pmos w=250u l=0.13u ng=25 m=1
.ends
.end
